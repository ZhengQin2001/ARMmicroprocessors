
module source_prob (
	probe);	

	input	[31:0]	probe;
endmodule
